`timescale 1ns/1ns
module astable_clock(output reg clk);
   
  initial clk = 0;
  always #5 clk = ~clk;

endmodule